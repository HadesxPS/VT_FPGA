//*****************************************************************************
// COPYRIGHT (c) 2013, Xiamen Tianma Microelectronics Co, Ltd
//
// File name     :  mux_decode.v
// Module name   :  mux_decode
//
// Author        :  sijian_luo
// Email         :  sijian_luo@tianma.cn
// Version       :  v 1.0
//
// Function      :  mux decoder
// Called by     :  --
//
// ----------------------------------------------------------------------------
// Revison
// 2014-08-01    :  create file
//*****************************************************************************
module mux_decode(
    input                 clk               ,
    input                 da                ,
    input                 db                ,
    output reg [1:0]      a
);

//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
// parameters
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++


//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
// variable declaration
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++


//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
// continuous assignment
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++


//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
// module instantiation
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++


//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
// block statement
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

//-----------------------------------------------------------------------------
// decoder
//-----------------------------------------------------------------------------
always @(posedge clk)
begin
    case ({da, db})
        2'b00:
        begin
            a <= 2'b01;
        end
        2'b01:
        begin
            a <= 2'b11;
        end
        2'b10:
        begin
            a <= 2'b10;
        end
        2'b11:
        begin
            a <= 2'b00;
        end
    endcase
end


endmodule