//*****************************************************************************
// COPYRIGHT (c) 2013, Xiamen Tianma Microelectronics Co, Ltd
//
// File name     :  clkrst.v
// Module name   :  clkrst
//
// Author        :  weipeng_wang
// Email         :  weipeng_wang@tianma.cn
// Version       :  v 1.0
//
// Function      :  clock and system reset generation
// Called by     :  --
//
// ----------------------------------------------------------------------------
// Revison
// 2015-06-17    :  create file
//*****************************************************************************
module clkrst (
    input                 clk_in            ,
    input                 rst_n_in          ,
    output                clk_sys           ,
    output reg            rst_n_sys
);

//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
// parameters
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
// variable declaration
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
reg                             rst_n_inclk                     ;
reg                             rst_n_sys_p1                    ;

//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
// continuous assignment
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
// module instantiation
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
mypll u_mypll(
    .inclk0                     ( clk_in                        ),
    .c0                         ( clk_sys                       )
);

//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
// block statement
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
always @(posedge clk_in)
begin
    rst_n_inclk <= rst_n_in;
end

always @(posedge clk_sys or negedge rst_n_inclk)
begin
    if (rst_n_inclk == 1'b0)
    begin
        rst_n_sys_p1 <= 1'b0;
        rst_n_sys    <= 1'b0;
    end
    else
    begin
        rst_n_sys_p1 <= 1'b1;
        rst_n_sys    <= rst_n_sys_p1;
    end
end

endmodule