library verilog;
use verilog.vl_types.all;
entity VT_Demo_vlg_tst is
end VT_Demo_vlg_tst;
